class packet extends uvm_sequence_item;

   `uvm_object_utils(packet)

endclass : packet
