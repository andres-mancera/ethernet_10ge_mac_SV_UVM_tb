`ifndef TEST_LIB__SVH
`define TEST_LIB__SVH

`include "../testcases/bringup_packet_test.sv"
`include "../testcases/oversized_packet_test.sv"
`include "../testcases/undersized_packet_test.sv"

`endif  // TEST_LIB__SVH
