`ifndef TEST_LIB__SVH
`define TEST_LIB__SVH

`include "../testcases/bringup_packet_test.sv"
`include "../testcases/oversized_packet_test.sv"
`include "../testcases/undersized_packet_test.sv"
`include "../testcases/small_large_packet_test.sv"
`include "../testcases/small_ipg_packet_test.sv"
`include "../testcases/zero_ipg_packet_test.sv"

`endif  // TEST_LIB__SVH
